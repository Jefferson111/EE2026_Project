`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.03.2019 20:54:05
// Design Name: 
// Module Name: Pause_Waveform
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Pause_Waveform(
    input [9:0] wave_sample,
    output reg [9:0] pause_sample = 0
    );
    
    
endmodule
